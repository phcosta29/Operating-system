module mux_controle_bios();
endmodule