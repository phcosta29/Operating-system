module mux_hd_bios();
endmodule