module memoriahd(input clk,
	input [9:0] setor_hd,
	input [15:0] endereco_hd,
	input [1:0] controle_hd,
	output [31:0] saida_instr
);
	reg[31:0]memoria[15:0][299:0];
	reg[15:0]endereco=16'b0000000000011111;	
	reg prim = 1'b0;

always@(posedge clk)
begin
	if(prim==1'b0)
	begin
		memoria[2][32]=32'b10101111110000000000000000001001; //loadi reg00001 valor=1 -> Verificado
		memoria[2][33]=32'b01110111110000000000000000001001; //print ula=1 -> Verificado
		memoria[2][34]=32'b10101111110000000000000000000110;
		memoria[2][35]=32'b01110111110000000000000000001010;	//loadi reg00010 valor=2 -> Verificado
		memoria[2][36]=32'b10101111110000000000000000001000; //load reg10000 valor=2 -> Verificado
		memoria[2][37]=32'b01110111110000000000000000001011; //print ula=2 -> Verificado
		memoria[2][38]=32'b10101111110000000000000000000111; //add reg00001+reg00010 valor=3 <- Verificado
		memoria[2][39]=32'b01110111110000000000000000001100; //print ula=3 -> Verificado 	
		memoria[2][40]=32'b10101111110000000000000000000100; //addi reg00011+1 valor=4 -> Verificado
		memoria[2][41]=32'b01110111110000000000000000000010; //print ula=4 -> Verificado
		memoria[2][42]=32'b01101111110000000000000000000010; //loadi reg00010 valor=1 -> Verificado
		memoria[2][43]=32'b00011000011111100000000000000001; //sub reg00011-reg00010 valor=3 <- Verificad
		memoria[2][44]=32'b01110000010000000000000000001000; //print ula=1 -> Verificado
		memoria[2][45]=32'b10101111110000000000000000000000; //sub reg00001-1 valor=2 <- Verificado
		memoria[2][46]=32'b01110111110000000000000000000011; //print ula=2 -> Verificado
		memoria[2][47]=32'b01101111110000000000000000000010; //jump pc0000000000010100 -> verificado
		memoria[2][48]=32'b00011000101111100000000000000010; //loadi reg00001 valor=1 -> Verificado
		memoria[2][49]=32'b01110000100000000000000000000111; //print ula=1 -> Verificado
		memoria[2][50]=32'b01101111000000000000000000000111; //loadi reg00001 valor=2 -> Verificado
		memoria[2][51]=32'b01101111110000000000000000000011; //loadi reg00010 valor=1 -> Verificado
		memoria[2][52]=32'b01011000111110011111000000000000; //and reg00010&reg00001 valor=0 -> Verificado
		memoria[2][53]=32'b10101111110000000000000000000001; //print ula=0 -> Verificado
		memoria[2][54]=32'b01001111110001100000000001010011; //andi reg00010&valor0000000000000001 valor=1 -> Verificado
		memoria[2][55]=32'b01101111000000000000000000000011; //print ula=1 -> Verificado	
		memoria[2][56]=32'b01110111000000000000000000000101; //or reg00010|reg00001 valor=3 -> Verificado
		memoria[2][57]=32'b01101111110000000000000000000011; //print ula=3 -> Verificado
		memoria[2][58]=32'b00001001001111100000000000000001; //ori reg00010|valor0000000000000001 valor=3 -> Verificado
		memoria[2][59]=32'b01110001000000000000000000000100; //print ula=3 -> Verificado
		memoria[2][60]=32'b01101111000000000000000000001000; //branch end0000000000101000 -> Verificado
		memoria[2][61]=32'b01101111110000000000000000000100; //branch not equal end0000000000101000 -> Verficado
		memoria[2][62]=32'b01011001011110011111000000000000; //loadi reg00001 valor=1 -> Verificado
		memoria[2][63]=32'b10101111110000000000000000000001; //print ula=1 -> Verificado
		memoria[2][64]=32'b01001111110010100000000000110100; //loadi reg00010 valor=2 -> Verificado
		memoria[2][65]=32'b10101111110000000000000000001001; //slt reg00001 e reg00010 valor=1 -> Verificado
		memoria[2][66]=32'b01101111100000000000000000000101; //print ula=1 -> Verificado
		memoria[2][67]=32'b00000111011111111110000000000000; //slti reg00001 valor0000000000000001 valor=0 -> Verificado
		memoria[2][68]=32'b11000111001110100000000000000000; //print ula=0 -> Verificado
		memoria[2][69]=32'b10101111110000000000000000001001; //not reg00001 valor=1 -> verificado
		memoria[2][70]=32'b01101111100000000000000000000100; //print ula=65534 -> Verificado
		memoria[2][71]=32'b00000111011111111110000000000000; //input valor=4
		memoria[2][72]=32'b11000111111110100000000000000000; //print ula=4 -> Verificado
		memoria[2][73]=32'b01011001101111111100000000000000;
		memoria[2][74]=32'b10101111110000000000000000000001;
		memoria[2][75]=32'b01001111110011000000000000101110;
		memoria[2][76]=32'b01000000000000000000000000110000;
		memoria[2][77]=32'b01101111000000000000000000000100;
		memoria[2][78]=32'b01110111000000000000000000000101;
		memoria[2][79]=32'b01101111110000000000000000000100;
		memoria[2][80]=32'b00001001111111100000000000000001;
		memoria[2][81]=32'b01110001110000000000000000000100;
		memoria[2][82]=32'b01000000000000000000000000011101;
		memoria[2][83]=32'b01101111000000000000000000000101;
		memoria[2][84]=32'b01101111110000000000000000000011;
		memoria[2][85]=32'b01001111111110000000000000111000;
		memoria[2][86]=32'b10101010000000000000000000000001;
		memoria[2][87]=32'b01000000000000000000000000111010;
		memoria[2][88]=32'b10101010000000000000000000000000;
		memoria[2][89]=32'b10101111110000000000000000000001;
		memoria[2][90]=32'b01001111110100000000000000111101;
		memoria[2][91]=32'b01000000000000000000000001001111;
		memoria[2][92]=32'b01101111110000000000000000000011;
		memoria[2][93]=32'b10101111100000000000000000001001;
		memoria[2][94]=32'b00000111011111111110000000000000;
		memoria[2][95]=32'b11000111001110100000000000000000;
		memoria[2][96]=32'b01110111000000000000000000000110;
		memoria[2][97]=32'b01101111110000000000000000000101;
		memoria[2][98]=32'b10101111100000000000000000001001;
		memoria[2][99]=32'b00000111011111111110000000000000;
		memoria[2][100]=32'b11000111001110100000000000000000;
		memoria[2][101]=32'b01101111110000000000000000000011;
		memoria[2][102]=32'b10101111100000000000000000001001;
		memoria[2][103]=32'b00000111011111111110000000000000;
		memoria[2][104]=32'b10000111001110100000000000000000;
		memoria[2][105]=32'b01101111000000000000000000000110;
		memoria[2][106]=32'b01101111110000000000000000000101;
		memoria[2][107]=32'b10101111100000000000000000001001;
		memoria[2][108]=32'b00000111011111111110000000000000;
		memoria[2][109]=32'b10000111001110100000000000000000;
		memoria[2][110]=32'b01101111110000000000000000000011;
		memoria[2][111]=32'b00001010011111100000000000000001;
		memoria[2][112]=32'b01110010010000000000000000000011;
		memoria[2][113]=32'b01000000000000000000000000010011;
		memoria[2][114]=32'b10001010110000000000000000000000;
		memoria[2][115]=32'b01110010110000000000000000001101;
		memoria[2][116]=32'b01101111110000000000000000001101;
		memoria[2][117]=32'b10101111100000000000000000001001;
		memoria[2][118]=32'b00000111011111111110000000000000;
		memoria[2][119]=32'b11000111001110100000000000000000;
		memoria[2][120]=32'b01110111000000000000000000001110;
		memoria[2][121]=32'b01101111110000000000000000001110;
		memoria[2][122]=32'b10010000001111100000000000000000;
		memoria[2][123]=32'b11111000000000000000000000000000;
		prim=1'b1;
	end
	if(controle_hd==2'b00)
		endereco=endereco+16'b0000000000000001;
	else
		endereco=16'b0000000000011111;
end
	assign saida_instr = memoria[setor_hd][endereco];
endmodule
